`timescale 1ns / 1ps

/*
Code for PS/2 Keyboard input obtained from:
http://www.instructables.com/id/PS2-Keyboard-for-FPGA/

Edited to fit TurfWars game controls.
*/

module keyboard(
    input CLOCK_50,
    input PS2_KBCLK,
    input PS2_KBDAT,
    output reg [4:0] KEY_PRESSED
   );

  // Specific Key codes
	wire [7:0] ARROW_UP = 8'h75;
	wire [7:0] ARROW_DOWN = 8'h72;
	wire [7:0] ARROW_LEFT = 8'h6B;
	wire [7:0] ARROW_RIGHT = 8'h74;
	wire [7:0] W = 8'h1D;
	wire [7:0] A = 8'h1C;
	wire [7:0] S = 8'h1B;
	wire [7:0] D = 8'h23;
	wire [7:0] Y = 8'h35;
	wire [7:0] G = 8'h34;
	wire [7:0] H = 8'h33;
	wire [7:0] J = 8'h3B;
	wire [7:0] P = 8'h4D;
	wire [7:0] L = 8'h4B;
	wire [7:0] COLON = 8'h4C;
	wire [7:0] QUOTES = 8'h52;
	wire [7:0] SPACE = 8'h29;

	reg read;				//this is 1 if still waits to receive more bits
	reg [11:0] count_reading;		//this is used to detect how much time passed since it received the previous codeword
	reg PREVIOUS_STATE;			//used to check the previous state of the keyboard clock signal to know if it changed
	reg scan_err;				//this becomes one if an error was received somewhere in the packet
	reg [10:0] scan_code;			//this stores 11 received bits
	reg [7:0] CODEWORD;			//this stores only the DATA codeword
	reg TRIG_ARR;				//this is triggered when full 11 bits are received
	reg [3:0]COUNT;				//tells how many bits were received until now (from 0 to 11)
	reg TRIGGER = 0;			//This acts as a 250 times slower than the board clock.
	reg [7:0]DOWNCOUNTER = 0;		//This is used together with TRIGGER - look the code

	//Set initial values
	initial begin
		PREVIOUS_STATE = 1;
		scan_err = 0;
		scan_code = 0;
		COUNT = 0;
		CODEWORD = 0;
		KEY_PRESSED = 0;
		read = 0;
		count_reading = 0;
	end

	always @(posedge CLOCK_50) begin				//This reduces the frequency 250 times
		if (DOWNCOUNTER < 249) begin			//and uses variable TRIGGER as the new board clock
			DOWNCOUNTER <= DOWNCOUNTER + 1;
			TRIGGER <= 0;
		end
		else begin
			DOWNCOUNTER <= 0;
			TRIGGER <= 1;
		end
	end

	always @(posedge CLOCK_50) begin
		if (TRIGGER) begin
			if (read)				//if it still waits to read full packet of 11 bits, then (read == 1)
				count_reading <= count_reading + 1;	//and it counts up this variable
			else 						//and later if check to see how big this value is.
				count_reading <= 0;			//if it is too big, then it resets the received data
		end
	end

	always @(posedge CLOCK_50) begin
	if (TRIGGER) begin						//If the down counter (CLK/250) is ready
		if (PS2_KBCLK != PREVIOUS_STATE) begin			//if the state of Clock pin changed from previous state
			if (!PS2_KBCLK) begin				//and if the keyboard clock is at falling edge
				read <= 1;				//mark down that it is still reading for the next bit
				scan_err <= 0;				//no errors
				scan_code[10:0] <= {PS2_KBDAT, scan_code[10:1]};	//add up the data received by shifting bits and adding one new bit
				COUNT <= COUNT + 1;			//
			end
		end
		else if (COUNT == 11) begin				//if it already received 11 bits
			COUNT <= 0;
			read <= 0;					//mark down that reading stopped
			TRIG_ARR <= 1;					//trigger out that the full pack of 11bits was received
			//calculate scan_err using parity bit
			if (!scan_code[10] || scan_code[0] || !(scan_code[1]^scan_code[2]^scan_code[3]^scan_code[4]
				^scan_code[5]^scan_code[6]^scan_code[7]^scan_code[8]
				^scan_code[9]))
				scan_err <= 1;
			else
				scan_err <= 0;
		end
		else  begin						//if it yet not received full pack of 11 bits
			TRIG_ARR <= 0;					//tell that the packet of 11bits was not received yet
			if (COUNT < 11 && count_reading >= 4000) begin	//and if after a certain time no more bits were received, then
				COUNT <= 0;				//reset the number of bits received
				read <= 0;				//and wait for the next packet
			end
		end
	PREVIOUS_STATE <= PS2_KBCLK;					//mark down the previous state of the keyboard clock
	end
	end

	always @(posedge CLOCK_50) begin
		if (TRIGGER) begin					//if the 250 times slower than board clock triggers
			if (TRIG_ARR) begin				//and if a full packet of 11 bits was received
				if (scan_err) begin			//BUT if the packet was NOT OK
					CODEWORD <= 8'd0;		//then reset the codeword register
				end
				else begin
					CODEWORD <= scan_code[8:1];	//else drop down the unnecessary  bits and transport the 7 DATA bits to CODEWORD reg
				end				//notice, that the codeword is also reversed! This is because the first bit to received
			end					//is supposed to be the last bit in the codeword…
			else CODEWORD <= 8'd0;				//not a full packet received, thus reset codeword
		end
		else CODEWORD <= 8'd0;					//no clock trigger, no data…
	end

  // Controls for TurfWars
	always @(posedge CLOCK_50) begin
		if (CODEWORD == ARROW_UP)
			KEY_PRESSED <= 5'd0;
		else if (CODEWORD == ARROW_DOWN)
			KEY_PRESSED <= 5'd1;
		else if (CODEWORD == ARROW_LEFT)
			KEY_PRESSED <= 5'd2;
		else if (CODEWORD == ARROW_RIGHT)
			KEY_PRESSED <= 5'd3;
		else if (CODEWORD == W)
			KEY_PRESSED <= 5'd4;
		else if (CODEWORD == S)
			KEY_PRESSED <= 5'd5;
		else if (CODEWORD == A)
			KEY_PRESSED <= 5'd6;
		else if (CODEWORD == D)
			KEY_PRESSED <= 5'd7;
		else if (CODEWORD == Y)
			KEY_PRESSED <= 5'd8;
		else if (CODEWORD == H)
			KEY_PRESSED <= 5'd9;
		else if (CODEWORD == G)
			KEY_PRESSED <= 5'd10;
		else if (CODEWORD == J)
			KEY_PRESSED <= 5'd11;
		else if (CODEWORD == P)
			KEY_PRESSED <= 5'd12;
		else if (CODEWORD == COLON)
			KEY_PRESSED <= 5'd13;
		else if (CODEWORD == L)
			KEY_PRESSED <= 5'd14;
		else if (CODEWORD == QUOTES)
			KEY_PRESSED <= 5'd15;
		else if (CODEWORD == SPACE)
			KEY_PRESSED <= 5'd16;
	end

endmodule
